interface intf(input logic clk, reset);
  logic [3:0] in1, in2;
  logic [4:0] out;
endinterface
