`include "sequence_item.sv"
`include "sequence1.sv"
`include "sequence2.sv"
`include "sequence3.sv"
`include "sequencer.sv"
`include "driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"
`include "agent.sv"
`include "environment.sv"
